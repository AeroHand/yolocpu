import lc3b_types::*;

module or_gate (output wire f, input wire a, b);

assign f = a || b;

endmodule : or_gate